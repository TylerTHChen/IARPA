module waves(
    input osc, // clock
    output logic GDS, // GDS Wave
    output logic QMOD, // QMOD Wave
    output logic clk
);

    logic reset;
    logic locked;
	
    clk_wiz_0 instance_name
   (
    // Clock out ports
    .clk(clk),     // output clk
    // Status and control signals
    .reset(reset), // input reset
    .locked(locked),       // output locked
   // Clock in ports
    .osc(osc)      // input osc
);
    // Define parameters for the size of waveforms and bit sequence
    parameter BIT = 823; 
    parameter WAVE = 8;

    // Sequence
    logic [WAVE-1:0] seq;
    assign seq = 8'b0101_0101;

    logic [0:BIT-1]bit0;
    logic [0:BIT-1]bit1;
    logic [0:BIT-1]QM;

/*
    // Initial block to load data from CSV files
    initial begin 
        $readmemb("GDS_0_50_d15_35_d10_30_d10_27_1.0u_100k.mem", bit0);
        $readmemb("GDS_1_50_d15_35_d10_30_d10_27_1.0u_100k.mem", bit1);
        $readmemb("Qmod_1.0u_100k_2498.mem",QM);
    end
*/

assign bit0 = 823'b1111000011110000111100001111000011110000111110001111100011110000111110001111100011110000111110001111100011110000111100001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign bit1 = 823'b0000111100001111000011110000111100001111100011110000111110001111000011111000111100001111100011110000111110001111000011110000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000001100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000011100000111000001110000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign QM = 823'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000;    // Counters
    integer bit_cnt = 0; 
    integer wave_cnt = 0;       

    // Always block to generate waveforms
    always @(posedge clk) begin
        if (bit_cnt < BIT) begin
            if (seq[wave_cnt] == 1'b1) begin
                GDS <= bit1[bit_cnt];
            end else begin
                GDS <= bit0[bit_cnt];
            end
            QMOD <= QM[bit_cnt];
            bit_cnt <= bit_cnt + 1;
            if (bit_cnt == BIT) begin
                bit_cnt <= 0;
                if(wave_cnt == WAVE)
                    wave_cnt <= 0;
                else
                    wave_cnt <= wave_cnt + 1;
            end
        end else begin
            // Reset counters when the sequence is complete
            bit_cnt <= 0;
            wave_cnt <= 0;
        end
    end
endmodule
